library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY cafeteira is
    Generic(
		a: INTEGER := 4	
    );
   Port ( 
		b : std_LOGIC
    );
	END cafeteira;
	
architecture behavioral of cafeteira is
	Begin
end behavioral;